`timescale 1ns / 1ps

module BranchUnit #(
    parameter PC_W = 9
) (
    input logic [PC_W-1:0] Cur_PC,
    input logic [31:0] Imm,
    input logic Branch,
    input logic jump,
    input logic jalrSel,
    input logic [31:0] AluResult,
    output logic [31:0] PC_Imm,
    output logic [31:0] PC_Four,
    output logic [31:0] BrPC,
    output logic PcSel
);

  logic Branch_Sel;
  logic [31:0] PC_Full;

  assign PC_Full = {23'b0, Cur_PC};
  assign PC_Imm = (jalrSel) ? (AluResult&(~(32'b001))) : (PC_Full + Imm);
  assign PC_Four = PC_Full + 32'b100;
  assign Branch_Sel = ((Branch && AluResult[0]) || (jump));

  assign BrPC = (Branch_Sel) ? PC_Imm : 32'b0;  // Branch -> PC+Imm   // Otherwise, BrPC value is not important
  assign PcSel = Branch_Sel;  // 1:branch is taken; 0:branch is not taken(choose pc+4)

  //assign PC_Imm = rs1 + IMM --> PC_Full = rs1; --> PC_Full = SrcA --> PC_Imm = AluResult;

endmodule
